module lab1(
  input wire 