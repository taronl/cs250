module asynchronous_reset(
  