
// demo1.v  My first project
// Author: Taron Linge & new comment
module demo1(
  input a,
  output reg y
);
  
  assign y = a;
  
endmodule