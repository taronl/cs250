module lab2(